// Generated build timestamp
`define BUILD_DATETIME "20250706153513"
